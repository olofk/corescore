`default_nettype none
module corescore_generic
(
 input wire  i_clk,
 input wire  i_rst,
 output wire o_uart_tx);

   parameter memfile_emitter = "emitter.hex";

   wire [7:0]  tdata;
   wire        tlast;
   wire        tvalid;
   wire        tready;

   corescorecore corescorecore
     (.i_clk     (i_clk),
      .i_rst     (i_rst),
      .o_tdata   (tdata),
      .o_tlast   (tlast),
      .o_tvalid  (tvalid),
      .i_tready  (tready));

   emitter_uart emitter
     (.i_clk     (i_clk),
      .i_rst     (i_rst),
      .i_tdata   (tdata),
      //.i_tlast   (tlast),
      .i_tvalid  (tvalid),
      .o_tready  (tready),
      .o_uart_tx (o_uart_tx));

endmodule
